module instruction_decode (read_data_1, read_data_2, extended_address,
 next_instruction, write_data);

output reg [31:0] read_data_1, read_data_2, extended_address;
input [31:0] next_instruction, write_data;


endmodule

