module instruction_fetch (next_instruction ,next_address, new_address);
//Starting


output reg [31:0] next_instruction, next_address;
input [31:0] new_address;


endmodule
