module execute (new_address, zero, alu_result, next_address,
 read_data_1, read_data_2, extended_address);

output reg [31:0] new_address, alu_result, next_address;
output reg zero; 
input [31:0] read_data_1, read_data_2, extended_address;



endmodule