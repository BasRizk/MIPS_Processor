module memory_access (read_data, new_address, zero, address_mem, write_data);

output reg [31:0] read_data;
input zero;
input [31:0] new_address, address_mem, write_data;



endmodule